/* CPU testbench */
`include "cpu.v"

module test;
    initial begin
        $display("Bad: cpu test not implemented");
    end
endmodule
