/* CPU testbench */
`include "cpu.v"
`include "alu.v"
`include "register.v"

module test;
    initial begin
        $display("Bad: cpu test not implemented");
    end
endmodule
